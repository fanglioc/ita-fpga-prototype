`timescale 1ns / 1ps

module expand_engine #(
    parameter INPUT_DIM = 64,
    parameter OUTPUT_DIM = 128,
    parameter WEIGHT_BITS = 4,
    parameter ACT_BITS = 8
)(
    input  logic clk,
    input  logic rst_n,
    input  logic [ACT_BITS-1:0] input_vec [INPUT_DIM],
    input  logic input_valid,
    output logic input_ready,
    output logic [ACT_BITS-1:0] output_vec [OUTPUT_DIM],
    output logic output_valid
);

    // State machine
    typedef enum logic [1:0] {
        IDLE,
        COMPUTE,
        DONE
    } state_t;
    
    state_t state;
    
    // Weight storage (Block RAM)
    // 128 neurons × 64 weights × 4 bits = 32 Kbits = 4 BRAM36
    logic [WEIGHT_BITS-1:0] weights [OUTPUT_DIM][INPUT_DIM];
    
    // Initialize weights from file (generated by Python)
    initial begin
        $readmemh("../weights/weights_expand.hex", weights);
    end
    
    // Computation counter
    logic [$clog2(INPUT_DIM):0] compute_cnt;
    
    // Parallel MAC units
    logic [ACT_BITS+WEIGHT_BITS+$clog2(INPUT_DIM)-1:0] accumulators [OUTPUT_DIM];
    logic [ACT_BITS+WEIGHT_BITS-1:0] mult_results [OUTPUT_DIM];
    
    // Generate MAC array
    genvar i;
    generate
        for (i = 0; i < OUTPUT_DIM; i++) begin : mac_array
            // Constant-coefficient multiplier
            assign mult_results[i] = input_vec[compute_cnt] * weights[i][compute_cnt];
            
            // Accumulator
            always_ff @(posedge clk) begin
                if (state == IDLE) begin
                    accumulators[i] <= 0;
                end else if (state == COMPUTE) begin
                    accumulators[i] <= accumulators[i] + mult_results[i];
                end
            end
            
            // Output with ReLU and saturation
            always_ff @(posedge clk) begin
                if (state == DONE) begin
                    if (accumulators[i][ACT_BITS+WEIGHT_BITS+$clog2(INPUT_DIM)-1]) begin
                        // Negative (sign bit set) → ReLU = 0
                        output_vec[i] <= 0;
                    end else begin
                        // Positive → saturate to ACT_BITS
                        logic [ACT_BITS+WEIGHT_BITS+$clog2(INPUT_DIM)-1:0] shifted;
                        shifted = accumulators[i] >> WEIGHT_BITS;  // Scale back
                        if (shifted > 255) begin
                            output_vec[i] <= 255;
                        end else begin
                            output_vec[i] <= shifted[ACT_BITS-1:0];
                        end
                    end
                end
            end
        end
    endgenerate
    
    // Control FSM
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            compute_cnt <= 0;
            output_valid <= 0;
        end else begin
            case (state)
                IDLE: begin
                    output_valid <= 0;
                    if (input_valid) begin
                        state <= COMPUTE;
                        compute_cnt <= 0;
                    end
                end
                
                COMPUTE: begin
                    compute_cnt <= compute_cnt + 1;
                    if (compute_cnt == INPUT_DIM - 1) begin
                        state <= DONE;
                    end
                end
                
                DONE: begin
                    output_valid <= 1;
                    state <= IDLE;
                end
            endcase
        end
    end
    
    assign input_ready = (state == IDLE);
    
endmodule
